// megafunction wizard: %40G/100G Ethernet Intel FPGA IP v19.1%
// GENERATION: XML
// fortygig_eth_mac.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module fortygig_eth_mac (
		input  wire         clk_ref,               //             clk_ref.clk
		input  wire         pma_arst_ST,           //         pma_arst_ST.pma_arst_ST
		input  wire         pcs_rx_arst_ST,        //      pcs_rx_arst_ST.pcs_rx_arst_ST
		input  wire         pcs_tx_arst_ST,        //      pcs_tx_arst_ST.pcs_tx_arst_ST
		output wire [367:0] reconfig_from_xcvr,    //  reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [559:0] reconfig_to_xcvr,      //    reconfig_to_xcvr.reconfig_to_xcvr
		input  wire         clk_status,            //              status.clk
		input  wire [15:0]  status_addr,           //                    .address
		input  wire         status_read,           //                    .read
		input  wire         status_write,          //                    .write
		input  wire [31:0]  status_writedata,      //                    .writedata
		output wire [31:0]  status_readdata,       //                    .readdata
		output wire         status_readdata_valid, //                    .readdatavalid
		output wire         rx_inc_runt,           //              rx_inc.rx_inc_runt
		output wire         rx_inc_64,             //                    .rx_inc_64
		output wire         rx_inc_127,            //                    .rx_inc_127
		output wire         rx_inc_255,            //                    .rx_inc_255
		output wire         rx_inc_511,            //                    .rx_inc_511
		output wire         rx_inc_1023,           //                    .rx_inc_1023
		output wire         rx_inc_1518,           //                    .rx_inc_1518
		output wire         rx_inc_max,            //                    .rx_inc_max
		output wire         rx_inc_over,           //                    .rx_inc_over
		output wire         rx_inc_mcast_data_err, //                    .rx_inc_mcast_data_err
		output wire         rx_inc_mcast_data_ok,  //                    .rx_inc_mcast_data_ok
		output wire         rx_inc_bcast_data_err, //                    .rx_inc_bcast_data_err
		output wire         rx_inc_bcast_data_ok,  //                    .rx_inc_bcast_data_ok
		output wire         rx_inc_ucast_data_err, //                    .rx_inc_ucast_data_err
		output wire         rx_inc_ucast_data_ok,  //                    .rx_inc_ucast_data_ok
		output wire         rx_inc_mcast_ctrl,     //                    .rx_inc_mcast_ctrl
		output wire         rx_inc_bcast_ctrl,     //                    .rx_inc_bcast_ctrl
		output wire         rx_inc_ucast_ctrl,     //                    .rx_inc_ucast_ctrl
		output wire         rx_inc_pause,          //                    .rx_inc_pause
		output wire         rx_inc_fcs_err,        //                    .rx_inc_fcs_err
		output wire         rx_inc_fragment,       //                    .rx_inc_fragment
		output wire         rx_inc_jabber,         //                    .rx_inc_jabber
		output wire         rx_inc_sizeok_fcserr,  //                    .rx_inc_sizeok_fcserr
		output wire         tx_inc_64,             //              tx_inc.tx_inc_64
		output wire         tx_inc_127,            //                    .tx_inc_127
		output wire         tx_inc_255,            //                    .tx_inc_255
		output wire         tx_inc_511,            //                    .tx_inc_511
		output wire         tx_inc_1023,           //                    .tx_inc_1023
		output wire         tx_inc_1518,           //                    .tx_inc_1518
		output wire         tx_inc_max,            //                    .tx_inc_max
		output wire         tx_inc_over,           //                    .tx_inc_over
		output wire         tx_inc_mcast_data_err, //                    .tx_inc_mcast_data_err
		output wire         tx_inc_mcast_data_ok,  //                    .tx_inc_mcast_data_ok
		output wire         tx_inc_bcast_data_err, //                    .tx_inc_bcast_data_err
		output wire         tx_inc_bcast_data_ok,  //                    .tx_inc_bcast_data_ok
		output wire         tx_inc_ucast_data_err, //                    .tx_inc_ucast_data_err
		output wire         tx_inc_ucast_data_ok,  //                    .tx_inc_ucast_data_ok
		output wire         tx_inc_mcast_ctrl,     //                    .tx_inc_mcast_ctrl
		output wire         tx_inc_bcast_ctrl,     //                    .tx_inc_bcast_ctrl
		output wire         tx_inc_ucast_ctrl,     //                    .tx_inc_ucast_ctrl
		output wire         tx_inc_pause,          //                    .tx_inc_pause
		output wire         tx_inc_fcs_err,        //                    .tx_inc_fcs_err
		output wire         tx_inc_fragment,       //                    .tx_inc_fragment
		output wire         tx_inc_jabber,         //                    .tx_inc_jabber
		output wire         tx_inc_sizeok_fcserr,  //                    .tx_inc_sizeok_fcserr
		input  wire         pause_insert_tx,       //               pause.pause_insert_tx
		input  wire [15:0]  pause_insert_time,     //                    .pause_insert_time
		input  wire         pause_insert_mcast,    //                    .pause_insert_mcast
		input  wire [47:0]  pause_insert_dst,      //                    .pause_insert_dst
		input  wire [47:0]  pause_insert_src,      //                    .pause_insert_src
		output wire         remote_fault_status,   // remote_fault_status.remote_fault_status
		output wire         local_fault_status,    //  local_fault_status.local_fault_status
		input  wire         clk_rxmac,             //           clk_rxmac.clk_rxmac
		input  wire         clk_txmac,             //           clk_txmac.clk_txmac
		input  wire         mac_rx_arst_ST,        //      mac_rx_arst_ST.mac_rx_arst_ST
		input  wire         mac_tx_arst_ST,        //      mac_tx_arst_ST.mac_tx_arst_ST
		output wire [255:0] l4_rx_data,            //               l4_rx.l4_rx_data
		output wire [4:0]   l4_rx_empty,           //                    .l4_rx_empty
		output wire         l4_rx_startofpacket,   //                    .l4_rx_startofpacket
		output wire         l4_rx_endofpacket,     //                    .l4_rx_endofpacket
		output wire         l4_rx_error,           //                    .l4_rx_error
		output wire         l4_rx_valid,           //                    .l4_rx_valid
		output wire         l4_rx_fcs_valid,       //                    .l4_rx_fcs_valid
		output wire         l4_rx_fcs_error,       //                    .l4_rx_fcs_error
		input  wire [255:0] l4_tx_data,            //               l4_tx.l4_tx_data
		input  wire [4:0]   l4_tx_empty,           //                    .l4_tx_empty
		input  wire         l4_tx_startofpacket,   //                    .l4_tx_startofpacket
		input  wire         l4_tx_endofpacket,     //                    .l4_tx_endofpacket
		output wire         l4_tx_ready,           //                    .l4_tx_ready
		input  wire         l4_tx_valid,           //                    .l4_tx_valid
		output wire [3:0]   tx_serial,             //           tx_serial.tx_serial
		input  wire [3:0]   rx_serial,             //           rx_serial.rx_serial
		output wire         lanes_deskewed,        //      lanes_deskewed.lanes_deskewed
		output wire         tx_lanes_stable        //     tx_lanes_stable.tx_lanes_stable
	);

	wire        fortygig_eth_mac_inst_tx_lanes_stable_phy; // port fragment
	wire        fortygig_eth_mac_inst_lanes_deskewed_phy;  // port fragment
	wire  [3:0] fortygig_eth_mac_inst_tx_serial_reg;       // port fragment

	alt_e40_top #(
		.DEVICE_FAMILY          ("Stratix V"),
		.VARIANT                (3),
		.PHY_PLL                ("ATX"),
		.REF_CLK_FREQ           ("644.53125 MHz"),
		.ENABLE_STATISTICS_CNTR (1),
		.en_synce_support       (0),
		.HAS_ADAPTERS           (1),
		.IS_CAUI4               (0),
		.TO_XCVR_WIDTH          (560),
		.FROM_XCVR_WIDTH        (368),
		.FAST_SIMULATION        (0),
		.STATUS_CLK_KHZ         (125000),
		.HAS_MAC                (1),
		.HAS_PHY                (1),
		.ENA_KR4                (0),
		.SYNTH_SEQ              (1),
		.SYNTH_FEC              (0),
		.SYNTH_AN               (1),
		.SYNTH_LT               (1),
		.LINK_TIMER_KR          (504),
		.OPTIONAL_RXEQ          (0),
		.BERWIDTH               (12),
		.TRNWTWIDTH             (7),
		.MAINTAPWIDTH           (6),
		.POSTTAPWIDTH           (5),
		.PRETAPWIDTH            (4),
		.VMAXRULE               (60),
		.VMINRULE               (9),
		.VODMINRULE             (24),
		.VPOSTRULE              (31),
		.VPRERULE               (15),
		.PREMAINVAL             (60),
		.PREPOSTVAL             (0),
		.PREPREVAL              (0),
		.INITMAINVAL            (52),
		.INITPOSTVAL            (30),
		.INITPREVAL             (5),
		.AN_CHAN                (1),
		.AN_PAUSE               (3),
		.AN_TECH                (8),
		.AN_FEC                 (0),
		.ERR_INDICATION         (1),
		.FEC_USE_M20K           (1)
	) fortygig_eth_mac_inst (
		.clk_ref                  (clk_ref),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //             clk_ref.clk
		.pma_arst_ST              (pma_arst_ST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         pma_arst_ST.pma_arst_ST
		.pcs_rx_arst_ST           (pcs_rx_arst_ST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //      pcs_rx_arst_ST.pcs_rx_arst_ST
		.pcs_tx_arst_ST           (pcs_tx_arst_ST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //      pcs_tx_arst_ST.pcs_tx_arst_ST
		.reconfig_from_xcvr       (reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //  reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr         (reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //    reconfig_to_xcvr.reconfig_to_xcvr
		.clk_status               (clk_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //              status.clk
		.status_addr              (status_addr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .address
		.status_read              (status_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .read
		.status_write             (status_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .write
		.status_writedata         (status_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                    .writedata
		.status_readdata          (status_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                    .readdata
		.status_readdata_valid    (status_readdata_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .readdatavalid
		.rx_inc_runt              (rx_inc_runt),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //              rx_inc.rx_inc_runt
		.rx_inc_64                (rx_inc_64),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .rx_inc_64
		.rx_inc_127               (rx_inc_127),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rx_inc_127
		.rx_inc_255               (rx_inc_255),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rx_inc_255
		.rx_inc_511               (rx_inc_511),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rx_inc_511
		.rx_inc_1023              (rx_inc_1023),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .rx_inc_1023
		.rx_inc_1518              (rx_inc_1518),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .rx_inc_1518
		.rx_inc_max               (rx_inc_max),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rx_inc_max
		.rx_inc_over              (rx_inc_over),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .rx_inc_over
		.rx_inc_mcast_data_err    (rx_inc_mcast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .rx_inc_mcast_data_err
		.rx_inc_mcast_data_ok     (rx_inc_mcast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .rx_inc_mcast_data_ok
		.rx_inc_bcast_data_err    (rx_inc_bcast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .rx_inc_bcast_data_err
		.rx_inc_bcast_data_ok     (rx_inc_bcast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .rx_inc_bcast_data_ok
		.rx_inc_ucast_data_err    (rx_inc_ucast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .rx_inc_ucast_data_err
		.rx_inc_ucast_data_ok     (rx_inc_ucast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .rx_inc_ucast_data_ok
		.rx_inc_mcast_ctrl        (rx_inc_mcast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .rx_inc_mcast_ctrl
		.rx_inc_bcast_ctrl        (rx_inc_bcast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .rx_inc_bcast_ctrl
		.rx_inc_ucast_ctrl        (rx_inc_ucast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .rx_inc_ucast_ctrl
		.rx_inc_pause             (rx_inc_pause),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .rx_inc_pause
		.rx_inc_fcs_err           (rx_inc_fcs_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .rx_inc_fcs_err
		.rx_inc_fragment          (rx_inc_fragment),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                    .rx_inc_fragment
		.rx_inc_jabber            (rx_inc_jabber),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .rx_inc_jabber
		.rx_inc_sizeok_fcserr     (rx_inc_sizeok_fcserr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .rx_inc_sizeok_fcserr
		.tx_inc_64                (tx_inc_64),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //              tx_inc.tx_inc_64
		.tx_inc_127               (tx_inc_127),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .tx_inc_127
		.tx_inc_255               (tx_inc_255),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .tx_inc_255
		.tx_inc_511               (tx_inc_511),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .tx_inc_511
		.tx_inc_1023              (tx_inc_1023),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .tx_inc_1023
		.tx_inc_1518              (tx_inc_1518),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .tx_inc_1518
		.tx_inc_max               (tx_inc_max),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .tx_inc_max
		.tx_inc_over              (tx_inc_over),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .tx_inc_over
		.tx_inc_mcast_data_err    (tx_inc_mcast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .tx_inc_mcast_data_err
		.tx_inc_mcast_data_ok     (tx_inc_mcast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .tx_inc_mcast_data_ok
		.tx_inc_bcast_data_err    (tx_inc_bcast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .tx_inc_bcast_data_err
		.tx_inc_bcast_data_ok     (tx_inc_bcast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .tx_inc_bcast_data_ok
		.tx_inc_ucast_data_err    (tx_inc_ucast_data_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .tx_inc_ucast_data_err
		.tx_inc_ucast_data_ok     (tx_inc_ucast_data_ok),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .tx_inc_ucast_data_ok
		.tx_inc_mcast_ctrl        (tx_inc_mcast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .tx_inc_mcast_ctrl
		.tx_inc_bcast_ctrl        (tx_inc_bcast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .tx_inc_bcast_ctrl
		.tx_inc_ucast_ctrl        (tx_inc_ucast_ctrl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .tx_inc_ucast_ctrl
		.tx_inc_pause             (tx_inc_pause),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .tx_inc_pause
		.tx_inc_fcs_err           (tx_inc_fcs_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .tx_inc_fcs_err
		.tx_inc_fragment          (tx_inc_fragment),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                    .tx_inc_fragment
		.tx_inc_jabber            (tx_inc_jabber),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .tx_inc_jabber
		.tx_inc_sizeok_fcserr     (tx_inc_sizeok_fcserr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .tx_inc_sizeok_fcserr
		.pause_insert_tx          (pause_insert_tx),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //               pause.pause_insert_tx
		.pause_insert_time        (pause_insert_time),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .pause_insert_time
		.pause_insert_mcast       (pause_insert_mcast),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                    .pause_insert_mcast
		.pause_insert_dst         (pause_insert_dst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                    .pause_insert_dst
		.pause_insert_src         (pause_insert_src),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                    .pause_insert_src
		.remote_fault_status      (remote_fault_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   // remote_fault_status.remote_fault_status
		.local_fault_status       (local_fault_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //  local_fault_status.local_fault_status
		.clk_rxmac                (clk_rxmac),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           clk_rxmac.clk_rxmac
		.clk_txmac                (clk_txmac),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           clk_txmac.clk_txmac
		.mac_rx_arst_ST           (mac_rx_arst_ST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //      mac_rx_arst_ST.mac_rx_arst_ST
		.mac_tx_arst_ST           (mac_tx_arst_ST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //      mac_tx_arst_ST.mac_tx_arst_ST
		.l4_rx_data               (l4_rx_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //               l4_rx.l4_rx_data
		.l4_rx_empty              (l4_rx_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_rx_empty
		.l4_rx_startofpacket      (l4_rx_startofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .l4_rx_startofpacket
		.l4_rx_endofpacket        (l4_rx_endofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .l4_rx_endofpacket
		.l4_rx_error              (l4_rx_error),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_rx_error
		.l4_rx_valid              (l4_rx_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_rx_valid
		.l4_rx_fcs_valid          (l4_rx_fcs_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                    .l4_rx_fcs_valid
		.l4_rx_fcs_error          (l4_rx_fcs_error),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                    .l4_rx_fcs_error
		.l4_tx_data               (l4_tx_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //               l4_tx.l4_tx_data
		.l4_tx_empty              (l4_tx_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_tx_empty
		.l4_tx_startofpacket      (l4_tx_startofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .l4_tx_startofpacket
		.l4_tx_endofpacket        (l4_tx_endofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .l4_tx_endofpacket
		.l4_tx_ready              (l4_tx_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_tx_ready
		.l4_tx_valid              (l4_tx_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .l4_tx_valid
		.tx_serial_reg            (fortygig_eth_mac_inst_tx_serial_reg[3:0]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //           tx_serial.tx_serial
		.rx_serial_reg            (rx_serial[3:0]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //           rx_serial.rx_serial
		.lanes_deskewed_phy       (fortygig_eth_mac_inst_lanes_deskewed_phy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //      lanes_deskewed.lanes_deskewed
		.tx_lanes_stable_phy      (fortygig_eth_mac_inst_tx_lanes_stable_phy),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //     tx_lanes_stable.tx_lanes_stable
		.rx_clk_ref               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_clk_ref               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.rx_recovered_clk         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.pll_locked               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_serial_clk            (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.reconfig_from_xcvr0      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.reconfig_to_xcvr0        (210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                               //         (terminated)
		.reconfig_from_xcvr1      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.reconfig_to_xcvr1        (210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                               //         (terminated)
		.reconfig_from_xcvr2      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.reconfig_to_xcvr2        (210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                               //         (terminated)
		.reconfig_from_xcvr3      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.reconfig_to_xcvr3        (210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                               //         (terminated)
		.pause_match_from_rx      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.pause_time_from_rx       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.remote_fault_from_rx     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.local_fault_from_rx      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.remote_fault_to_tx       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.local_fault_to_tx        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.pause_match_to_tx        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.pause_time_to_tx         (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.rx_mii_valid_mac         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.rx_mii_valid_phy         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.rx_mii_d_mac             (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                 //         (terminated)
		.rx_mii_d_phy             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.rx_mii_c_mac             (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.rx_mii_c_phy             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.lanes_deskewed_mac       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_mii_d_phy             (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                 //         (terminated)
		.tx_mii_d_mac             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.tx_mii_c_phy             (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_mii_c_mac             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.tx_mii_valid_phy         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_mii_valid_mac         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.tx_mii_ready_mac         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.tx_mii_ready_phy         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.tx_lanes_stable_mac      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.l8_rx_data               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_empty              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_startofpacket      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_endofpacket        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_error              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_valid              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_fcs_valid          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_rx_fcs_error          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_tx_data               (512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.l8_tx_empty              (6'b000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //         (terminated)
		.l8_tx_startofpacket      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.l8_tx_endofpacket        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.l8_tx_ready              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.l8_tx_valid              (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.din                      (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                 //         (terminated)
		.din_start                (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //         (terminated)
		.din_end_pos              (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.din_ack                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_d                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_c                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_first_data          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_last_data           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_runt_last_data      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_payload             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_fcs_error           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_fcs_valid           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_dst_addr_match      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dout_valid               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.a10_reconfig_write       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.a10_reconfig_read        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.a10_reconfig_address     (12'b000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.a10_reconfig_writedata   (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.a10_reconfig_readdata    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.a10_reconfig_waitrequest (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.rc_busy                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.lt_start_rc              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.main_rc                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.post_rc                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.pre_rc                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.tap_to_upd               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.en_lcl_rxeq              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.rxeq_done                (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.seq_start_rc             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.pcs_mode_rc              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.reco_mif_done            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //         (terminated)
		.upi_mode_en              (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_adj                  (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.upi_inc                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_dec                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_pre                  (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_init                 (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_st_bert              (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_train_err            (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_lock_err             (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upi_rx_trained           (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         (terminated)
		.upo_enable               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_frame_lock           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_cm_done              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_bert_done            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_ber_cnt              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_ber_max              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.upo_coef_max             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dfe_start_rc             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.dfe_mode                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.ctle_start_rc            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.ctle_rc                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //         (terminated)
		.ctle_mode                ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //         (terminated)
	);

	assign tx_lanes_stable = { fortygig_eth_mac_inst_tx_lanes_stable_phy };

	assign lanes_deskewed = { fortygig_eth_mac_inst_lanes_deskewed_phy };

	assign tx_serial = { fortygig_eth_mac_inst_tx_serial_reg[3:0] };

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2021 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="alt_e40_e100" version="19.1" >
// Retrieval info: 	<generic name="DEVICE_FAMILY" value="Stratix V" />
// Retrieval info: 	<generic name="MAC_CONFIG" value="40 Gbe" />
// Retrieval info: 	<generic name="CORE_OPTION" value="MAC &amp; PHY" />
// Retrieval info: 	<generic name="PHY_CONFIG" value="1" />
// Retrieval info: 	<generic name="INTERFACE" value="Avalon-ST Interface" />
// Retrieval info: 	<generic name="VARIANT" value="3" />
// Retrieval info: 	<generic name="PHY_PLL" value="ATX" />
// Retrieval info: 	<generic name="PHY_REFCLK" value="1" />
// Retrieval info: 	<generic name="STATUS_CLK_KHZ_SIV" value="50.0" />
// Retrieval info: 	<generic name="STATUS_CLK_KHZ_SV" value="125.0" />
// Retrieval info: 	<generic name="ENABLE_STATISTICS_CNTR" value="1" />
// Retrieval info: 	<generic name="en_synce_support" value="0" />
// Retrieval info: 	<generic name="ENA_KR4_gui" value="0" />
// Retrieval info: 	<generic name="SYNTH_SEQ" value="1" />
// Retrieval info: 	<generic name="SYNTH_FEC" value="0" />
// Retrieval info: 	<generic name="SYNTH_AN_gui" value="1" />
// Retrieval info: 	<generic name="SYNTH_LT_gui" value="1" />
// Retrieval info: 	<generic name="LINK_TIMER_KR" value="504" />
// Retrieval info: 	<generic name="OPTIONAL_UP" value="0" />
// Retrieval info: 	<generic name="OPTIONAL_RXEQ" value="0" />
// Retrieval info: 	<generic name="BERWIDTH_gui" value="4095" />
// Retrieval info: 	<generic name="TRNWTWIDTH_gui" value="127" />
// Retrieval info: 	<generic name="MAINTAPWIDTH" value="6" />
// Retrieval info: 	<generic name="POSTTAPWIDTH" value="5" />
// Retrieval info: 	<generic name="PRETAPWIDTH" value="4" />
// Retrieval info: 	<generic name="VMAXRULE" value="60" />
// Retrieval info: 	<generic name="VMINRULE" value="9" />
// Retrieval info: 	<generic name="VODMINRULE" value="24" />
// Retrieval info: 	<generic name="VPOSTRULE" value="31" />
// Retrieval info: 	<generic name="VPRERULE" value="15" />
// Retrieval info: 	<generic name="PREMAINVAL" value="60" />
// Retrieval info: 	<generic name="PREPOSTVAL" value="0" />
// Retrieval info: 	<generic name="PREPREVAL" value="0" />
// Retrieval info: 	<generic name="INITMAINVAL" value="52" />
// Retrieval info: 	<generic name="INITPOSTVAL" value="30" />
// Retrieval info: 	<generic name="INITPREVAL" value="5" />
// Retrieval info: 	<generic name="AN_GIGE" value="0" />
// Retrieval info: 	<generic name="AN_XAUI" value="0" />
// Retrieval info: 	<generic name="AN_BASER" value="0" />
// Retrieval info: 	<generic name="AN_40GBP" value="1" />
// Retrieval info: 	<generic name="AN_40GCR" value="0" />
// Retrieval info: 	<generic name="AN_100G" value="0" />
// Retrieval info: 	<generic name="AN_CHAN" value="1" />
// Retrieval info: 	<generic name="AN_PAUSE_C0" value="1" />
// Retrieval info: 	<generic name="AN_PAUSE_C1" value="1" />
// Retrieval info: 	<generic name="AN_SELECTOR" value="1" />
// Retrieval info: 	<generic name="CAPABLE_FEC" value="1" />
// Retrieval info: 	<generic name="ENABLE_FEC" value="1" />
// Retrieval info: 	<generic name="ERR_INDICATION" value="1" />
// Retrieval info: 	<generic name="FEC_USE_M20K" value="1" />
// Retrieval info: </instance>
// IPFS_FILES : fortygig_eth_mac.vo
// RELATED_FILES: fortygig_eth_mac.v, alt_e40_top.v, alt_e40_bridge.v, alt_e40_lock_timer.v, alt_e40_status_sync.v, alt_e40_sticky_flag.v, alt_e40_sync_arst.v, alt_e40_user_mode_det.v, alt_e40_adapter_rx.v, alt_e40_wide_l4if_rx2to4.v, alt_e40_wide_l4if_rx2to4fifo.v, alt_e40_wide_l4if_rxfifo.v, alt_e40_wide_l4if_sopfifo.v, alt_e40_adapter_tx.v, alt_e40_wide_l4if_tx4to2.v, alt_e40_wide_l4if_tx4to2fifo.v, alt_e40_wide_l4if_txfifo.v, alt_e40_mac.v, alt_e40_crc32_d64_sig.v, alt_e40_crc32_rev_1.v, alt_e40_crc32_rev_2.v, alt_e40_crc32_rev_4.v, alt_e40_crc32_z64_x1.v, alt_e40_crc32_z64_x2.v, alt_e40_fcs_40g.v, alt_e40_insert_parity.v, alt_e40_mlab_delay.v, alt_e40_mlab_sr_cells.v, alt_e40_remove_parity.v, alt_e40_reverse_words.v, alt_e40_six_three_comp.v, alt_e40_stat_cntr_1port.v, alt_e40_stat_cntr_2port.v, alt_e40_mac_addr_regs.v, alt_e40_mac_csr.v, alt_e40_status_cntr_pause_sync.v, alt_e40_doe_cmd_fifo.v, alt_e40_doe_fifo.v, alt_e40_doe_storage_ram.v, alt_e40_dst_addr_chk.v, alt_e40_m9k_with_par.v, alt_e40_mac_link_fault_det.v, alt_e40_mac_link_fault_det_ns.v, alt_e40_mac_rx.v, alt_e40_mac_rx_stats.v, alt_e40_pause_chk.v, alt_e40_runt_comparator.v, alt_e40_runt_detect.v, alt_e40_rx_inspect_40g.v, alt_e40_rx_pad_strip.v, alt_e40_rx_preamble_passthrough.v, alt_e40_gap_monitor.v, alt_e40_gap_monitor_ns.v, alt_e40_idle_count.v, alt_e40_mac_link_fault_gen.v, alt_e40_mac_tx.v, alt_e40_mac_tx_stats.v, alt_e40_pause_dp.v, alt_e40_pause_ebuf.v, alt_e40_sum_of_3bit_pair.v, alt_e40_twelve_four_comp.v, alt_e40_tx_pad_and_spacer.v, alt_e40_tx_preamble_passthrough.v, alt_e40_tx_to_mii.v, alt_e40_xlgmii_rom.v, alt_e40_phy_pma_sv.v, alt_e40_pma_sv_bridge.v, alt_e40_phy.v, alt_e40_frequency_monitor.v, alt_e40_phy_csr.v, alt_e40_status_cntr_sync.v, alt_e40_sticky_flag_group.v, alt_e40_phy_pcs.v, alt_e40_gray_to_bin.v, alt_e40_mlab_dcfifo.v, alt_e40_mlab_fifo_cells.v, alt_e40_random_delay.v, alt_e40_block_decoder.v, alt_e40_block_decoder_ns.v, alt_e40_descrambler.v, alt_e40_framed_descrambler.v, alt_e40_gearbox_40_66.v, alt_e40_lane_marker_compare.v, alt_e40_lane_marker_lock.v, alt_e40_mii_decode_multiple.v, alt_e40_pcs_ber.v, alt_e40_pcs_ber_cnt_ns.v, alt_e40_pcs_ber_sm.v, alt_e40_pcs_rx.v, alt_e40_pcs_rx_testmode.v, alt_e40_prbs_rx.v, alt_e40_reorder_destripe.v, alt_e40_rx_lane.v, alt_e40_rx_lane_array.v, alt_e40_rx_nav_region.v, alt_e40_word_align_control.v, alt_e40_block_encoder.v, alt_e40_block_encoder_ns.v, alt_e40_framed_scrambler.v, alt_e40_gearbox_66_40.v, alt_e40_mii_encode_multiple.v, alt_e40_pcs_tx.v, alt_e40_prbs_tx.v, alt_e40_scrambler.v, alt_e40_tx_lane.v, alt_e40_tx_lane_array.v, alt_e40_tx_nav_region.v, alt_e40_e4x10.v, altera_xcvr_functions.sv, altera_xcvr_low_latency_phy.sv, alt_pma_controller_tgx.v, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, sv_xcvr_low_latency_phy_nr.sv, sv_xcvr_10g_custom_native.sv, sv_xcvr_custom_native.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
